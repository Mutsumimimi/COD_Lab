`define PDU_IMEM_FILE "D:\code_field\COD_Lab\Lab3\PDU_v3-main\vsrc\inits\pdu_inits\riscv\pdu_imem.ini"
`define PDU_DMEM_FILE "D:\code_field\COD_Lab\Lab3\PDU_v3-main\vsrc\inits\pdu_inits\riscv\pdu_dmem.ini"
`define CPU_IMEM_FILE "D:\code_field\COD_Lab\Lab3\PDU_v3-main\vsrc\inits\cpu_inits\instr.ini"
`define CPU_DMEM_FILE "D:\code_field\COD_Lab\Lab3\PDU_v3-main\vsrc\inits\cpu_inits\data.ini"